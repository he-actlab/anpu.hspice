**** Design of a Resistor Network ****
.subckt ResNetwork8b   Iout_resDAC     dacIin   w0in    w1in   w2in  w3in  w4in  w5in  w6in  w7in
r0    dacIin    net2240    res_ntwk
r1    net2240   net2241    res_ntwk
r2    net2241   net2242    res_ntwk
r3    net2242   net2243    res_ntwk
r4    net2243   net2244    res_ntwk
r5    net2244   net2245    res_ntwk
r6    net2245   net2246    res_ntwk
r7    net2246   net2247    res_ntwk
r8    net2247   net2248    res_ntwk
r9    net2248   net2249    res_ntwk
r10    net2249   net2250    res_ntwk
r11    net2250   net2251    res_ntwk
r12    net2251   net2252    res_ntwk
r13    net2252   net2253    res_ntwk
r14    net2253   net2254    res_ntwk
r15    net2254   net2255    res_ntwk
r16    net2255   net2256    res_ntwk
r17    net2256   net2257    res_ntwk
r18    net2257   net2258    res_ntwk
r19    net2258   net2259    res_ntwk
r20    net2259   net2260    res_ntwk
r21    net2260   net2261    res_ntwk
r22    net2261   net2262    res_ntwk
r23    net2262   net2263    res_ntwk
r24    net2263   net2264    res_ntwk
r25    net2264   net2265    res_ntwk
r26    net2265   net2266    res_ntwk
r27    net2266   net2267    res_ntwk
r28    net2267   net2268    res_ntwk
r29    net2268   net2269    res_ntwk
r30    net2269   net2270    res_ntwk
r31    net2270   net2271    res_ntwk
r32    net2271   net2272    res_ntwk
r33    net2272   net2273    res_ntwk
r34    net2273   net2274    res_ntwk
r35    net2274   net2275    res_ntwk
r36    net2275   net2276    res_ntwk
r37    net2276   net2277    res_ntwk
r38    net2277   net2278    res_ntwk
r39    net2278   net2279    res_ntwk
r40    net2279   net2280    res_ntwk
r41    net2280   net2281    res_ntwk
r42    net2281   net2282    res_ntwk
r43    net2282   net2283    res_ntwk
r44    net2283   net2284    res_ntwk
r45    net2284   net2285    res_ntwk
r46    net2285   net2286    res_ntwk
r47    net2286   net2287    res_ntwk
r48    net2287   net2288    res_ntwk
r49    net2288   net2289    res_ntwk
r50    net2289   net2290    res_ntwk
r51    net2290   net2291    res_ntwk
r52    net2291   net2292    res_ntwk
r53    net2292   net2293    res_ntwk
r54    net2293   net2294    res_ntwk
r55    net2294   net2295    res_ntwk
r56    net2295   net2296    res_ntwk
r57    net2296   net2297    res_ntwk
r58    net2297   net2298    res_ntwk
r59    net2298   net2299    res_ntwk
r60    net2299   net2300    res_ntwk
r61    net2300   net2301    res_ntwk
r62    net2301   net2302    res_ntwk
r63    net2302   net2303    res_ntwk
r64    net2303   net2304    res_ntwk
r65    net2304   net2305    res_ntwk
r66    net2305   net2306    res_ntwk
r67    net2306   net2307    res_ntwk
r68    net2307   net2308    res_ntwk
r69    net2308   net2309    res_ntwk
r70    net2309   net2310    res_ntwk
r71    net2310   net2311    res_ntwk
r72    net2311   net2312    res_ntwk
r73    net2312   net2313    res_ntwk
r74    net2313   net2314    res_ntwk
r75    net2314   net2315    res_ntwk
r76    net2315   net2316    res_ntwk
r77    net2316   net2317    res_ntwk
r78    net2317   net2318    res_ntwk
r79    net2318   net2319    res_ntwk
r80    net2319   net2320    res_ntwk
r81    net2320   net2321    res_ntwk
r82    net2321   net2322    res_ntwk
r83    net2322   net2323    res_ntwk
r84    net2323   net2324    res_ntwk
r85    net2324   net2325    res_ntwk
r86    net2325   net2326    res_ntwk
r87    net2326   net2327    res_ntwk
r88    net2327   net2328    res_ntwk
r89    net2328   net2329    res_ntwk
r90    net2329   net2310    res_ntwk
r91    net2330   net2331    res_ntwk
r92    net2331   net2332    res_ntwk
r93    net2332   net2333    res_ntwk
r94    net2333   net2334    res_ntwk
r95    net2334   net2335    res_ntwk
r96    net2335   net2336    res_ntwk
r97    net2336   net2337    res_ntwk
r98    net2337   net2338    res_ntwk
r99    net2338   net2339    res_ntwk
r100   net2339   net2340    res_ntwk
r101   net2340   net2341    res_ntwk
r102   net2341   net2342    res_ntwk
r103   net2342   net2343    res_ntwk
r104   net2343   net2344    res_ntwk
r105   net2344   net2345    res_ntwk
r106   net2345   net2346    res_ntwk
r107   net2346   net2347    res_ntwk
r108   net2347   net2348    res_ntwk
r109   net2348   net2349    res_ntwk
r110   net2349   net2350    res_ntwk
r111   net2350   net2351    res_ntwk
r112   net2351   net2352    res_ntwk
r113   net2352   net2353    res_ntwk
r114   net2353   net2354    res_ntwk
r115   net2354   net2355    res_ntwk
r116   net2355   net2356    res_ntwk
r117   net2356   net2357    res_ntwk
r118   net2357   net2358    res_ntwk
r119   net2358   net2359    res_ntwk
r120   net2359   net2360    res_ntwk
r121   net2360   net2361    res_ntwk
r122   net2361   net2362    res_ntwk
r123   net2362   net2363    res_ntwk
r124   net2363   net2364    res_ntwk
r125   net2364   net2365    res_ntwk
r126   net2365   net2366    res_ntwk
r127   net2366   net2367    res_ntwk
r128   net2367   net2368    res_ntwk
r129   net2368   net2369    res_ntwk
r130   net2369   net2370    res_ntwk
r131   net2370   net2371    res_ntwk
r132   net2371   net2372    res_ntwk
r133   net2372   net2373    res_ntwk
r134   net2373   net2374    res_ntwk
r135   net2374   net2375    res_ntwk
r136   net2375   net2376    res_ntwk
r137   net2376   net2377    res_ntwk
r138   net2377   net2378    res_ntwk
r139   net2378   net2379    res_ntwk
r140   net2379   net2380    res_ntwk
r141   net2380   net2381    res_ntwk
r142   net2481   net2382    res_ntwk
r143   net2482   net2383    res_ntwk
r144   net2483   net2384    res_ntwk
r145   net2484   net2385    res_ntwk
r146   net2485   net2386    res_ntwk
r147   net2486   net2387    res_ntwk
r148   net2487   net2388    res_ntwk
r149   net2488   net2389    res_ntwk
r150   net2389   net2390    res_ntwk
r151   net2390   net2391    res_ntwk
r152   net2391   net2392    res_ntwk
r153   net2392   net2393    res_ntwk
r154   net2393   net2394    res_ntwk
r155   net2394   net2395    res_ntwk
r156   net2395   net2396    res_ntwk
r157   net2396   net2397    res_ntwk
r158   net2397   net2398    res_ntwk
r159   net2398   net2399    res_ntwk
r160   net2399   net2400    res_ntwk
r161   net2400   net2401    res_ntwk
r162   net2401   net2402    res_ntwk
r163   net2402   net2403    res_ntwk
r164   net2403   net2404    res_ntwk
r165   net2404   net2405    res_ntwk
r166   net2405   net2406    res_ntwk
r167   net2406   net2407    res_ntwk
r168   net2407   net2408    res_ntwk
r169   net2408   net2409    res_ntwk
r170   net2409   net2410    res_ntwk
r171   net2410   net2411    res_ntwk
r172   net2411   net2412    res_ntwk
r173   net2412   net2413    res_ntwk
r174   net2413   net2414    res_ntwk
r175   net2414   net2415    res_ntwk
r176   net2415   net2416    res_ntwk
r177   net2416   net2417    res_ntwk
r178   net2417   net2418    res_ntwk
r179   net2418   net2419    res_ntwk
r180   net2419   net2420    res_ntwk
r181   net2420   net2421    res_ntwk
r182   net2421   net2422    res_ntwk
r183   net2422   net2423    res_ntwk
r184   net2423   net2424    res_ntwk
r185   net2424   net2425    res_ntwk
r186   net2425   net2426    res_ntwk
r187   net2426   net2427    res_ntwk
r188   net2427   net2428    res_ntwk
r189   net2428   net2429    res_ntwk
r190   net2429   net2430    res_ntwk
r191   net2430   net2431    res_ntwk
r192   net2431   net2432    res_ntwk
r193   net2432   net2433    res_ntwk
r194   net2433   net2434    res_ntwk
r195   net2434   net2435    res_ntwk
r196   net2435   net2436    res_ntwk
r197   net2436   net2437    res_ntwk
r198   net2437   net2438    res_ntwk
r199   net2438   net2439    res_ntwk
r200   net2439   net2440    res_ntwk
r201   net2440   net2441    res_ntwk
r202   net2441   net2442    res_ntwk
r203   net2442   net2443    res_ntwk
r204   net2443   net2444    res_ntwk
r205   net2444   net2445    res_ntwk
r206   net2445   net2446    res_ntwk
r207   net2446   net2447    res_ntwk
r208   net2447   net2448    res_ntwk
r209   net2448   net2449    res_ntwk
r210   net2449   net2450    res_ntwk
r211   net2450   net2451    res_ntwk
r212   net2451   net2452    res_ntwk
r213   net2452   net2453    res_ntwk
r214   net2453   net2454    res_ntwk
r215   net2454   net2455    res_ntwk
r216   net2455   net2456    res_ntwk
r217   net2456   net2457    res_ntwk
r218   net2457   net2458    res_ntwk
r219   net2458   net2459    res_ntwk
r220   net2459   net2460    res_ntwk
r221   net2460   net2461    res_ntwk
r222   net2461   net2462    res_ntwk
r223   net2462   net2463    res_ntwk
r224   net2463   net2464    res_ntwk
r225   net2464   net2465    res_ntwk
r226   net2465   net2466    res_ntwk
r227   net2466   net2467    res_ntwk
r228   net2467   net2468    res_ntwk
r229   net2468   net2469    res_ntwk
r230   net2469   net2470    res_ntwk
r231   net2470   net2471    res_ntwk
r232   net2471   net2472    res_ntwk
r233   net2472   net2473    res_ntwk
r234   net2473   net2474    res_ntwk
r235   net2474   net2475    res_ntwk
r236   net2475   net2476    res_ntwk
r237   net2476   net2477    res_ntwk
r238   net2477   net2478    res_ntwk
r239   net2478   net2479    res_ntwk
r240   net2479   net2480    res_ntwk
r241   net2480   net2481    res_ntwk
r242   net2481   net2482    res_ntwk
r243   net2482   net2483    res_ntwk
r244   net2483   net2484    res_ntwk
r245   net2484   net2485    res_ntwk
r246   net2485   net2486    res_ntwk
r247   net2486   net2487    res_ntwk
r248   net2487   net2488    res_ntwk
r249   net2488   net2489    res_ntwk
r250   net2489   net2490    res_ntwk
r251   net2490   net2491    res_ntwk
r252   net2491   net2492    res_ntwk
r253   net2492   net2493    res_ntwk
r254   net2493   net2494    res_ntwk
r255   net2494   net2495    res_ntwk
v0     net2495   0          dc=Vbias_diffpair
I0     net2496   net2240    w0in   net2241    TxSwitch1to2_2
I1     net2497   net2242    w0in   net2243    TxSwitch1to2_2
I2     net2498   net2244    w0in   net2245    TxSwitch1to2_2
I3     net2499   net2246    w0in   net2247    TxSwitch1to2_2
I4     net2500   net2248    w0in   net2249    TxSwitch1to2_2
I5     net2501   net2250    w0in   net2251    TxSwitch1to2_2
I6     net2502   net2252    w0in   net2253    TxSwitch1to2_2
I7     net2503   net2254    w0in   net2255    TxSwitch1to2_2
I8     net2504   net2256    w0in   net2257    TxSwitch1to2_2
I9     net2505   net2258    w0in   net2259    TxSwitch1to2_2
I10    net2506   net2260    w0in   net2261    TxSwitch1to2_2
I11    net2507   net2262    w0in   net2263    TxSwitch1to2_2
I12    net2508   net2264    w0in   net2265    TxSwitch1to2_2
I13    net2509   net2266    w0in   net2267    TxSwitch1to2_2
I14    net2500   net2268    w0in   net2269    TxSwitch1to2_2
I15    net2511   net2270    w0in   net2271    TxSwitch1to2_2
I16    net2512   net2272    w0in   net2273    TxSwitch1to2_2
I17    net2513   net2274    w0in   net2275    TxSwitch1to2_2
I18    net2514   net2276    w0in   net2277    TxSwitch1to2_2
I19    net2515   net2278    w0in   net2279    TxSwitch1to2_2
I20    net2516   net2280    w0in   net2281    TxSwitch1to2_2
I21    net2517   net2282    w0in   net2283    TxSwitch1to2_2
I22    net2518   net2284    w0in   net2285    TxSwitch1to2_2
I23    net2519   net2286    w0in   net2287    TxSwitch1to2_2
I24    net2520   net2288    w0in   net2289    TxSwitch1to2_2
I25    net2521   net2290    w0in   net2291    TxSwitch1to2_2
I26    net2522   net2292    w0in   net2293    TxSwitch1to2_2
I27    net2523   net2294    w0in   net2295    TxSwitch1to2_2
I28    net2524   net2296    w0in   net2297    TxSwitch1to2_2
I29    net2525   net2298    w0in   net2299    TxSwitch1to2_2
I30    net2526   net2300    w0in   net2301    TxSwitch1to2_2
I31    net2527   net2302    w0in   net2303    TxSwitch1to2_2
I32    net2528   net2304    w0in   net2305    TxSwitch1to2_2
I33    net2529   net2306    w0in   net2307    TxSwitch1to2_2
I34    net2520   net2308    w0in   net2309    TxSwitch1to2_2
I35    net2531   net2310    w0in   net2311    TxSwitch1to2_2
I36    net2532   net2312    w0in   net2313    TxSwitch1to2_2
I37    net2533   net2314    w0in   net2315    TxSwitch1to2_2
I38    net2534   net2316    w0in   net2317    TxSwitch1to2_2
I39    net2535   net2318    w0in   net2319    TxSwitch1to2_2
I40    net2536   net2320    w0in   net2321    TxSwitch1to2_2
I41    net2537   net2322    w0in   net2323    TxSwitch1to2_2
I42    net2538   net2324    w0in   net2325    TxSwitch1to2_2
I43    net2539   net2326    w0in   net2327    TxSwitch1to2_2
I44    net2530   net2328    w0in   net2329    TxSwitch1to2_2
I45    net2541   net2330    w0in   net2331    TxSwitch1to2_2
I46    net2542   net2332    w0in   net2333    TxSwitch1to2_2
I47    net2543   net2334    w0in   net2335    TxSwitch1to2_2
I48    net2544   net2336    w0in   net2337    TxSwitch1to2_2
I49    net2545   net2338    w0in   net2339    TxSwitch1to2_2
I50    net2546   net2340    w0in   net2341    TxSwitch1to2_2
I51    net2547   net2342    w0in   net2343    TxSwitch1to2_2
I52    net2548   net2344    w0in   net2345    TxSwitch1to2_2
I53    net2549   net2346    w0in   net2347    TxSwitch1to2_2
I54    net2550   net2348    w0in   net2349    TxSwitch1to2_2
I55    net2551   net2350    w0in   net2351    TxSwitch1to2_2
I56    net2552   net2352    w0in   net2353    TxSwitch1to2_2
I57    net2553   net2354    w0in   net2355    TxSwitch1to2_2
I58    net2554   net2356    w0in   net2357    TxSwitch1to2_2
I59    net2555   net2358    w0in   net2359    TxSwitch1to2_2
I60    net2556   net2360    w0in   net2361    TxSwitch1to2_2
I61    net2557   net2362    w0in   net2363    TxSwitch1to2_2
I62    net2558   net2364    w0in   net2365    TxSwitch1to2_2
I63    net2559   net2366    w0in   net2367    TxSwitch1to2_2
I64    net2560   net2368    w0in   net2369    TxSwitch1to2_2
I65    net2561   net2370    w0in   net2371    TxSwitch1to2_2
I66    net2562   net2372    w0in   net2373    TxSwitch1to2_2
I67    net2563   net2374    w0in   net2375    TxSwitch1to2_2
I68    net2564   net2376    w0in   net2377    TxSwitch1to2_2
I69    net2565   net2378    w0in   net2379    TxSwitch1to2_2
I70    net2566   net2380    w0in   net2381    TxSwitch1to2_2
I71    net2567   net2382    w0in   net2383    TxSwitch1to2_2
I72    net2568   net2384    w0in   net2385    TxSwitch1to2_2
I73    net2569   net2386    w0in   net2387    TxSwitch1to2_2
I74    net2570   net2388    w0in   net2389    TxSwitch1to2_2
I75    net2571   net2390    w0in   net2391    TxSwitch1to2_2
I76    net2572   net2392    w0in   net2393    TxSwitch1to2_2
I77    net2573   net2394    w0in   net2395    TxSwitch1to2_2
I78    net2574   net2396    w0in   net2397    TxSwitch1to2_2
I79    net2575   net2398    w0in   net2399    TxSwitch1to2_2
I80    net2576   net2400    w0in   net2401    TxSwitch1to2_2
I81    net2577   net2402    w0in   net2403    TxSwitch1to2_2
I82    net2578   net2404    w0in   net2405    TxSwitch1to2_2
I83    net2579   net2406    w0in   net2407    TxSwitch1to2_2
I84    net2580   net2408    w0in   net2409    TxSwitch1to2_2
I85    net2581   net2410    w0in   net2411    TxSwitch1to2_2
I86    net2582   net2412    w0in   net2413    TxSwitch1to2_2
I87    net2583   net2414    w0in   net2415    TxSwitch1to2_2
I88    net2584   net2416    w0in   net2417    TxSwitch1to2_2
I89    net2585   net2418    w0in   net2419    TxSwitch1to2_2
I90    net2586   net2420    w0in   net2421    TxSwitch1to2_2
I91    net2587   net2422    w0in   net2423    TxSwitch1to2_2
I92    net2588   net2424    w0in   net2425    TxSwitch1to2_2
I93    net2589   net2426    w0in   net2427    TxSwitch1to2_2
I94    net2590   net2428    w0in   net2429    TxSwitch1to2_2
I95    net2591   net2430    w0in   net2431    TxSwitch1to2_2
I96    net2592   net2432    w0in   net2433    TxSwitch1to2_2
I97    net2593   net2434    w0in   net2435    TxSwitch1to2_2
I98    net2594   net2436    w0in   net2437    TxSwitch1to2_2
I99    net2595   net2438    w0in   net2439    TxSwitch1to2_2
I100   net2596   net2440    w0in   net2441    TxSwitch1to2_2
I101   net2597   net2442    w0in   net2443    TxSwitch1to2_2
I102   net2598   net2444    w0in   net2445    TxSwitch1to2_2
I103   net2599   net2446    w0in   net2447    TxSwitch1to2_2
I104   net2600   net2448    w0in   net2449    TxSwitch1to2_2
I105   net2601   net2450    w0in   net2451    TxSwitch1to2_2
I106   net2602   net2452    w0in   net2453    TxSwitch1to2_2
I107   net2603   net2454    w0in   net2455    TxSwitch1to2_2
I108   net2604   net2456    w0in   net2457    TxSwitch1to2_2
I109   net2605   net2458    w0in   net2459    TxSwitch1to2_2
I110   net2606   net2460    w0in   net2461    TxSwitch1to2_2
I111   net2607   net2462    w0in   net2463    TxSwitch1to2_2
I112   net2608   net2464    w0in   net2465    TxSwitch1to2_2
I113   net2609   net2466    w0in   net2467    TxSwitch1to2_2
I114   net2610   net2468    w0in   net2469    TxSwitch1to2_2
I115   net2611   net2470    w0in   net2471    TxSwitch1to2_2
I116   net2612   net2472    w0in   net2473    TxSwitch1to2_2
I117   net2613   net2474    w0in   net2475    TxSwitch1to2_2
I118   net2614   net2476    w0in   net2477    TxSwitch1to2_2
I119   net2615   net2478    w0in   net2479    TxSwitch1to2_2
I120    net2616   net2480    w0in   net2481    TxSwitch1to2_2
I121    net2617   net2482    w0in   net2483    TxSwitch1to2_2
I122    net2618   net2484    w0in   net2485    TxSwitch1to2_2
I123    net2619   net2486    w0in   net2487    TxSwitch1to2_2
I124    net2620   net2488    w0in   net2489    TxSwitch1to2_2
I125    net2621   net2490    w0in   net2491    TxSwitch1to2_2
I126    net2622   net2492    w0in   net2493    TxSwitch1to2_2
I127    net2623   net2494    w0in   net2495    TxSwitch1to2_2
I128    net2624   net2496    w0in   net2497    TxSwitch1to2_2
I129    net2625   net2498    w0in   net2499    TxSwitch1to2_2
I130    net2626   net2500    w0in   net2501    TxSwitch1to2_2
I131    net2627   net2502    w0in   net2503    TxSwitch1to2_2
I132    net2628   net2504    w0in   net2505    TxSwitch1to2_2
I133    net2629   net2506    w0in   net2507    TxSwitch1to2_2
I134    net2620   net2508    w0in   net2509    TxSwitch1to2_2
I135    net2631   net2510    w0in   net2511    TxSwitch1to2_2
I136    net2632   net2512    w0in   net2513    TxSwitch1to2_2
I137    net2633   net2514    w0in   net2515    TxSwitch1to2_2
I138    net2634   net2516    w0in   net2517    TxSwitch1to2_2
I139    net2635   net2518    w0in   net2519    TxSwitch1to2_2
I140    net2636   net2520    w0in   net2521    TxSwitch1to2_2
I141    net2637   net2522    w0in   net2523    TxSwitch1to2_2
I142    net2638   net2524    w0in   net2525    TxSwitch1to2_2
I143    net2639   net2526    w0in   net2527    TxSwitch1to2_2
I144    net2630   net2528    w0in   net2529    TxSwitch1to2_2
I145    net2641   net2530    w0in   net2531    TxSwitch1to2_2
I146    net2642   net2532    w0in   net2533    TxSwitch1to2_2
I147    net2643   net2534    w0in   net2535    TxSwitch1to2_2
I148    net2644   net2536    w0in   net2537    TxSwitch1to2_2
I149    net2645   net2538    w0in   net2539    TxSwitch1to2_2
I150    net2646   net2540    w0in   net2541    TxSwitch1to2_2
I151    net2647   net2542    w0in   net2543    TxSwitch1to2_2
I152    net2648   net2544    w0in   net2545    TxSwitch1to2_2
I153    net2649   net2546    w0in   net2547    TxSwitch1to2_2
I154    net2650   net2548    w0in   net2549    TxSwitch1to2_2
I155    net2651   net2550    w0in   net2551    TxSwitch1to2_2
I156    net2652   net2552    w0in   net2553    TxSwitch1to2_2
I157    net2653   net2554    w0in   net2555    TxSwitch1to2_2
I158    net2654   net2556    w0in   net2557    TxSwitch1to2_2
I159    net2655   net2558    w0in   net2559    TxSwitch1to2_2
I160    net2656   net2560    w0in   net2561    TxSwitch1to2_2
I161    net2657   net2562    w0in   net2563    TxSwitch1to2_2
I162    net2658   net2564    w0in   net2565    TxSwitch1to2_2
I163    net2659   net2566    w0in   net2567    TxSwitch1to2_2
I164    net2660   net2568    w0in   net2569    TxSwitch1to2_2
I165    net2661   net2570    w0in   net2571    TxSwitch1to2_2
I166    net2662   net2572    w0in   net2573    TxSwitch1to2_2
I167    net2663   net2574    w0in   net2575    TxSwitch1to2_2
I168    net2664   net2576    w0in   net2577    TxSwitch1to2_2
I169    net2665   net2578    w0in   net2579    TxSwitch1to2_2
I170    net2666   net2580    w0in   net2581    TxSwitch1to2_2
I171    net2667   net2582    w0in   net2583    TxSwitch1to2_2
I172    net2668   net2584    w0in   net2585    TxSwitch1to2_2
I173    net2669   net2586    w0in   net2587    TxSwitch1to2_2
I174    net2670   net2588    w0in   net2589    TxSwitch1to2_2
I175    net2671   net2590    w0in   net2591    TxSwitch1to2_2
I176    net2672   net2592    w0in   net2593    TxSwitch1to2_2
I177    net2673   net2594    w0in   net2595    TxSwitch1to2_2
I178    net2674   net2596    w0in   net2597    TxSwitch1to2_2
I179    net2675   net2598    w0in   net2599    TxSwitch1to2_2
I180    net2676   net2600    w0in   net2601    TxSwitch1to2_2
I181    net2677   net2602    w0in   net2603    TxSwitch1to2_2
I182    net2678   net2604    w0in   net2605    TxSwitch1to2_2
I183    net2679   net2606    w0in   net2607    TxSwitch1to2_2
I184    net2680   net2608    w0in   net2609    TxSwitch1to2_2
I185    net2681   net2610    w0in   net2611    TxSwitch1to2_2
I186    net2682   net2612    w0in   net2613    TxSwitch1to2_2
I187    net2683   net2614    w0in   net2615    TxSwitch1to2_2
I188    net2684   net2616    w0in   net2617    TxSwitch1to2_2
I189    net2685   net2618    w0in   net2619    TxSwitch1to2_2
I190    net2686   net2620    w0in   net2621    TxSwitch1to2_2
I191    net2687   net2622    w0in   net2623    TxSwitch1to2_2
I192    net2688   net2624    w0in   net2625    TxSwitch1to2_2
I193    net2689   net2626    w0in   net2627    TxSwitch1to2_2
I194    net2690   net2628    w0in   net2629    TxSwitch1to2_2
I195    net2691   net2630    w0in   net2631    TxSwitch1to2_2
I196    net2692   net2632    w0in   net2633    TxSwitch1to2_2
I197    net2693   net2634    w0in   net2635    TxSwitch1to2_2
I198    net2694   net2636    w0in   net2637    TxSwitch1to2_2
I199    net2695   net2638    w0in   net2639    TxSwitch1to2_2
I200   net2696   net2640    w0in   net2641    TxSwitch1to2_2
I201   net2697   net2642    w0in   net2643    TxSwitch1to2_2
I202   net2698   net2644    w0in   net2645    TxSwitch1to2_2
I203   net2699   net2646    w0in   net2647    TxSwitch1to2_2
I204   net2700   net2648    w0in   net2649    TxSwitch1to2_2
I205   net2701   net2650    w0in   net2651    TxSwitch1to2_2
I206   net2702   net2652    w0in   net2653    TxSwitch1to2_2
I207   net2703   net2654    w0in   net2655    TxSwitch1to2_2
I208   net2704   net2656    w0in   net2657    TxSwitch1to2_2
I209   net2705   net2658    w0in   net2659    TxSwitch1to2_2
I210   net2706   net2660    w0in   net2661    TxSwitch1to2_2
I211   net2707   net2662    w0in   net2663    TxSwitch1to2_2
I212   net2708   net2664    w0in   net2665    TxSwitch1to2_2
I213   net2709   net2666    w0in   net2667    TxSwitch1to2_2
I214   net2710   net2668    w0in   net2669    TxSwitch1to2_2
I215   net2711   net2670    w0in   net2671    TxSwitch1to2_2
I216   net2712   net2672    w0in   net2673    TxSwitch1to2_2
I217   net2713   net2674    w0in   net2675    TxSwitch1to2_2
I218   net2714   net2676    w0in   net2677    TxSwitch1to2_2
I219   net2715   net2678    w0in   net2679    TxSwitch1to2_2
I220   net2716   net2680    w0in   net2681    TxSwitch1to2_2
I221   net2717   net2682    w0in   net2683    TxSwitch1to2_2
I222   net2718   net2684    w0in   net2685    TxSwitch1to2_2
I223   net2719   net2686    w0in   net2687    TxSwitch1to2_2
I224   net2720   net2688    w0in   net2689    TxSwitch1to2_2
I225   net2721   net2690    w0in   net2691    TxSwitch1to2_2
I226   net2722   net2692    w0in   net2693    TxSwitch1to2_2
I227   net2723   net2694    w0in   net2695    TxSwitch1to2_2
I228   net2724   net2696    w0in   net2697    TxSwitch1to2_2
I229   net2725   net2698    w0in   net2699    TxSwitch1to2_2
I230   net2726   net2700    w0in   net2701    TxSwitch1to2_2
I231   net2727   net2702    w0in   net2703    TxSwitch1to2_2
I232   net2728   net2704    w0in   net2705    TxSwitch1to2_2
I233   net2729   net2706    w0in   net2707    TxSwitch1to2_2
I234   net2720   net2708    w0in   net2709    TxSwitch1to2_2
I235   net2731   net2710    w0in   net2711    TxSwitch1to2_2
I236   net2732   net2712    w0in   net2713    TxSwitch1to2_2
I237   net2733   net2714    w0in   net2715    TxSwitch1to2_2
I238   net2734   net2716    w0in   net2717    TxSwitch1to2_2
I239   net2735   net2718    w0in   net2719    TxSwitch1to2_2
I240   net2736   net2720    w0in   net2721    TxSwitch1to2_2
I241   net2737   net2722    w0in   net2723    TxSwitch1to2_2
I242   net2738   net2724    w0in   net2725    TxSwitch1to2_2
I243   net2739   net2726    w0in   net2727    TxSwitch1to2_2
I244   net2730   net2728    w0in   net2729    TxSwitch1to2_2
I245   net2741   net2730    w0in   net2731    TxSwitch1to2_2
I246   net2742   net2732    w0in   net2733    TxSwitch1to2_2
I247   net2743   net2734    w0in   net2735    TxSwitch1to2_2
I248   net2744   net2736    w0in   net2737    TxSwitch1to2_2
I249   net2745   net2738    w0in   net2739    TxSwitch1to2_2
I250   net2746   net2740    w0in   net2741    TxSwitch1to2_2
I251   net2747   net2742    w0in   net2743    TxSwitch1to2_2
I252   net2748   net2744    w0in   net2745    TxSwitch1to2_2
I253   net2749   net2746    w0in   net2747    TxSwitch1to2_2
I254   net2750   net2748    w0in   net2749    TxSwitch1to2_2
.ends ResNetwork8b