.subckt FlashADC6b_Vsrc_comp Vin_ADC fv_pos0	fv_pos1		fv_pos2		fv_pos3		fv_pos4		fv_pos5		fv_pos6
+									 fv_pos7 	fv_pos8		fv_pos9		fv_pos10	fv_pos11	fv_pos12	fv_pos13
+									 fv_pos14	fv_pos15	fv_pos16 	fv_pos17 	fv_pos18 	fv_pos19	fv_pos20
+									 fv_pos21 	fv_pos22 	fv_pos23 	fv_pos24 	fv_pos25 	fV_pos26 	fv_pos27
+									 fv_pos28 	fv_pos29 	fv_pos30 	fv_pos31 	fv_pos32 	fv_pos33 	fv_pos34
+ 									 fv_pos35 	fv_pos36 	fv_pos37 	fV_pos38 	fV_pos38 	fv_pos39 	fv_pos40
+									 fv_pos41	fv_pos42	fv_pos43	fv_pos44 	fv_pos45	fv_pos46	fv_pos47
+									 fv_pos48 	fv_pos49	fv_pos50	fv_pos51	fv_pos52	fv_pos53	fv_pos54
+									 fv_pos55 	fv_pos56	fv_pos57 	fv_pos58	fv_pos59 	fv_pos60 	fv_pos61
+									 net3200
+									 fv_neg0	fv_neg1		fv_neg2		fv_neg3		fv_neg4		fv_neg5		fv_neg6
+									 fv_neg7 	fv_neg8		fv_neg9		fv_neg10	fv_neg11	fv_neg12	fv_neg13
+									 fv_neg14	fv_neg15	fv_neg16 	fv_neg17 	fv_neg18 	fv_neg19	fv_neg20
+									 fv_neg21 	fv_neg22 	fv_neg23 	fv_neg24 	fv_neg25 	fV_neg26 	fv_neg27
+									 fv_neg28 	fv_neg29 	fv_neg30 	fv_neg31 	fv_neg32 	fv_neg33 	fv_neg34
+ 									 fv_neg35 	fv_neg36 	fv_neg37 	fV_neg38 	fV_neg38 	fv_neg39 	fv_neg40
+									 fv_neg41	fv_neg42	fv_neg43	fv_neg44 	fv_neg45	fv_neg46	fv_neg47
+									 fv_neg48 	fv_neg49	fv_neg50	fv_neg51	fv_neg52	fv_neg53	fv_neg54
+									 fv_neg55 	fv_neg56	fv_neg57 	fv_neg58	fv_neg59 	fv_neg60 	fv_neg61
+									 net3201    Vltch_In


I122		Vin_ADC 		Vref16		Vltch_In	fv_pos16 	fv_neg16	Comparator
I121		Vin_ADC 		Vref17		Vltch_In	fv_pos17 	fv_neg17	Comparator
I200		Vin_ADC 		net0636		Vltch_In	net3200 	net3201		Comparator
I127 		Vin_ADC			net348   	Vltch_In	fV_pos61    fv_neg61    Comparator
I128 		Vin_ADC         net0635		Vltch_In	fv_pos60	fv_neg60	Comparator
I129 		Vin_ADC         net346		Vltch_In	fv_pos59	fv_neg59	Comparator
I130 		Vin_ADC         net342		Vltch_In	fv_pos58	fv_neg58	Comparator
I131 		Vin_ADC         net340		Vltch_In	fv_pos57	fv_neg57	Comparator
I132 		Vin_ADC         net338		Vltch_In	fv_pos56	fv_neg56	Comparator
I133 		Vin_ADC         net360		Vltch_In	fv_pos55	fv_neg55	Comparator
I134 		Vin_ADC         net358		Vltch_In	fv_pos54	fv_neg54	Comparator
I135 		Vin_ADC         net356		Vltch_In	fv_pos53	fv_neg53	Comparator
I136 		Vin_ADC         net354		Vltch_In	fv_pos52	fv_neg52	Comparator
I137 		Vin_ADC         net352		Vltch_In	fv_pos51	fv_neg51	Comparator
I138 		Vin_ADC         net350		Vltch_In	fv_pos50	fv_neg50	Comparator
I101 		Vin_ADC         Vref18		Vltch_In	fv_pos18	fv_neg18	Comparator
I100 		Vin_ADC         Vref19		Vltch_In	fv_pos19	fv_neg19	Comparator
I99 		Vin_ADC         Vref20		Vltch_In	fv_pos20	fv_neg20	Comparator
I98 		Vin_ADC         Vref21		Vltch_In	fv_pos21	fv_neg21	Comparator
I97 		Vin_ADC         Vref22		Vltch_In	fv_pos22	fv_neg22	Comparator
I96 		Vin_ADC         Vref23		Vltch_In	fv_pos23	fv_neg23	Comparator
I76 		Vin_ADC         Vref24		Vltch_In	fv_pos24	fv_neg24	Comparator
I75 		Vin_ADC         Vref25		Vltch_In	fv_pos25	fv_neg25	Comparator
I74 		Vin_ADC         Vref26		Vltch_In	fv_pos26	fv_neg26	Comparator
I73 		Vin_ADC         Vref27		Vltch_In	fv_pos27	fv_neg27	Comparator
I72 		Vin_ADC         Vref28		Vltch_In	fv_pos28	fv_neg28	Comparator
I71 		Vin_ADC         Vref29		Vltch_In	fv_pos29	fv_neg29	Comparator
I67			Vin_ADC         Vref30		Vltch_In	fv_pos30	fv_neg30	Comparator
I66 		Vin_ADC         Vref15		Vltch_In	fv_pos15	fv_neg15	Comparator
I59 		Vin_ADC         Vref14		Vltch_In	fv_pos14	fv_neg14	Comparator
I58	 		Vin_ADC         Vref13		Vltch_In	fv_pos13	fv_neg13	Comparator
I51 		Vin_ADC         Vref12		Vltch_In	fv_pos12	fv_neg12	Comparator
I50 		Vin_ADC         Vref11		Vltch_In	fv_pos11	fv_neg11	Comparator
I43 		Vin_ADC         Vref10		Vltch_In	fv_pos10	fv_neg10	Comparator
I42 		Vin_ADC         Vref9		Vltch_In	fv_pos9 	fv_neg9 	Comparator
I35 		Vin_ADC         Vref8		Vltch_In	fv_pos8 	fv_neg8 	Comparator
I33 		Vin_ADC         Vref7		Vltch_In	fv_pos7 	fv_neg7 	Comparator
I25 		Vin_ADC         Vref6		Vltch_In	fv_pos6 	fv_neg6 	Comparator
I22 		Vin_ADC         Vref5		Vltch_In	fv_pos5 	fv_neg5 	Comparator
I156 		Vin_ADC         net330		Vltch_In	fv_pos42 	fv_neg42 	Comparator
I157 		Vin_ADC         net328		Vltch_In	fv_pos43 	fv_neg43 	Comparator
I158 		Vin_ADC         net326		Vltch_In	fv_pos44 	fv_neg44 	Comparator
I159 		Vin_ADC         net302		Vltch_In	fv_pos45 	fv_neg45 	Comparator
I160 		Vin_ADC         net300		Vltch_In	fv_pos46 	fv_neg46 	Comparator
I194 		Vin_ADC         net322		Vltch_In	fv_pos33 	fv_neg33 	Comparator
I162		Vin_ADC         net320		Vltch_In	fv_pos34 	fv_neg34 	Comparator
I163 		Vin_ADC         net318		Vltch_In	fv_pos32 	fv_neg32 	Comparator
I164 		Vin_ADC         net314		Vltch_In	fv_pos35 	fv_neg35 	Comparator
I165 		Vin_ADC         net312		Vltch_In	fv_pos36 	fv_neg36 	Comparator
I17 		Vin_ADC         Vref4 		Vltch_In 	fv_pos4 	fv_neg4 	Comparator
I166 		Vin_ADC 		net310 		Vltch_In 	fv_pos37 	fv_neg37  	Comparator
I167 		Vin_ADC 		net308 		Vltch_In 	fv_pos38 	fv_neg38  	Comparator
I168 		Vin_ADC 		net336 		Vltch_In 	fv_pos39 	fv_neg39  	Comparator
I169 		Vin_ADC 		net334 		Vltch_In 	fv_pos40 	fv_neg40  	Comparator
I170 		Vin_ADC 		net332 		Vltch_In 	fv_pos41 	fv_neg41  	Comparator
I171 		Vin_ADC 		net324 		Vltch_In 	fv_pos49 	fv_neg49  	Comparator
I172 		Vin_ADC 		net306 		Vltch_In 	fv_pos48 	fv_neg48  	Comparator
I173 		Vin_ADC 		net304 		Vltch_In 	fv_pos47 	fv_neg47  	Comparator
I174 		Vin_ADC 		net316 		Vltch_In 	fv_pos31 	fv_neg31  	Comparator
I5 			Vin_ADC 		Vref1 		Vltch_In 	fv_pos1  	fv_neg1  	Comparator
I193 		Vin_ADC 		Vref0 		Vltch_In 	fv_pos0  	fv_neg0  	Comparator
I13 		Vin_ADC 		Vref3 		Vltch_In 	fv_pos3  	fv_neg3  	Comparator
I9  		Vin_ADC 		Vref2 		Vltch_In 	fv_pos2  	fv_neg2  	Comparator
V32			net360 			0